module main

import buffer
import buffer.gap
import buffer.rope

fn main() {
	println('Hello World!')
}
