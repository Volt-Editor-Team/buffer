module gap

import math

pub fn (mut g GapBuffer) remove(cursor int, count int) {
	byte_index := g.char_to_byte_index(cursor)
	g.shift_gap_to(byte_index)
	total_bytes := g.to_string()[cursor..cursor + count].bytes().len
	g.gap.end = math.min(total_bytes, g.data.len)
}
